-- NNFFPGA_Network_secondModel_statics.vhd
-- This is an automatically generated file containing the constants for the neural network
-- The constants are generated form a Keras Network Object via the Network-2-FPGA.py script

-- Autor: Christian Woznik
-- E-Mail: christian.woznik@posteo.de
-- This file war created on 2021-12-01
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library work;
use work.NNFPGA_pkg.all;
use work.NNFPGA_statics.all;

package NNFFPGA_Network_secondModel_statics is
	-- Layer Informations
	constant c_networksecondModelLayerInformation : t_networkInformation(0 to 1) := (
			0 => (activationFunction => 1, inputCount => 63, neuronCount =>5),
			1 => (activationFunction => 3, inputCount => 5, neuronCount =>6));


	-- Weights Array
	constant c_networksecondModelWeights : t_variableSizeIntegerArray(0 to 355) := (
			--Layer 1
			--Neuron 1
			0 => -6,
			1 => 15,
			2 => 0,
			3 => 0,
			4 => -17,
			5 => -2,
			6 => -5,
			7 => -9,
			8 => 9,
			9 => 4,
			10 => 1,
			11 => 0,
			12 => -4,
			13 => -1,
			14 => -6,
			15 => 3,
			16 => -3,
			17 => -1,
			18 => 2,
			19 => 3,
			20 => -8,
			21 => -1,
			22 => 5,
			23 => 2,
			24 => -2,
			25 => 5,
			26 => 3,
			27 => -7,
			28 => -11,
			29 => -8,
			30 => 5,
			31 => -1,
			32 => -2,
			33 => -1,
			34 => -2,
			35 => -8,
			36 => 2,
			37 => 5,
			38 => 3,
			39 => 0,
			40 => 0,
			41 => -9,
			42 => 7,
			43 => 5,
			44 => -3,
			45 => 0,
			46 => -1,
			47 => -1,
			48 => -4,
			49 => -3,
			50 => -1,
			51 => -6,
			52 => -23,
			53 => 22,
			54 => -4,
			55 => -2,
			56 => -1,
			57 => 3,
			58 => 3,
			59 => 1,
			60 => 0,
			61 => -1,
			62 => -2,
			63 => 1,
			--Neuron 2
			64 => 9,
			65 => 1,
			66 => 3,
			67 => 10,
			68 => -5,
			69 => 8,
			70 => 4,
			71 => -5,
			72 => 6,
			73 => -6,
			74 => -4,
			75 => -7,
			76 => 8,
			77 => -4,
			78 => -3,
			79 => 3,
			80 => -4,
			81 => -3,
			82 => 10,
			83 => 6,
			84 => 5,
			85 => 6,
			86 => 1,
			87 => 8,
			88 => 2,
			89 => 3,
			90 => -7,
			91 => -9,
			92 => 2,
			93 => -3,
			94 => 2,
			95 => -2,
			96 => 6,
			97 => 1,
			98 => -3,
			99 => 0,
			100 => 7,
			101 => -5,
			102 => 9,
			103 => 6,
			104 => -2,
			105 => -7,
			106 => -1,
			107 => -3,
			108 => 5,
			109 => 9,
			110 => 7,
			111 => -7,
			112 => 6,
			113 => 9,
			114 => -4,
			115 => -3,
			116 => -3,
			117 => -2,
			118 => -7,
			119 => 6,
			120 => 9,
			121 => 5,
			122 => -1,
			123 => 5,
			124 => 6,
			125 => 7,
			126 => 7,
			127 => -2,
			--Neuron 3
			128 => 6,
			129 => -15,
			130 => 7,
			131 => 2,
			132 => 17,
			133 => 0,
			134 => 0,
			135 => -2,
			136 => 1,
			137 => -1,
			138 => 0,
			139 => 2,
			140 => -1,
			141 => 2,
			142 => -2,
			143 => 10,
			144 => 10,
			145 => -2,
			146 => -4,
			147 => -5,
			148 => -12,
			149 => 4,
			150 => -5,
			151 => 5,
			152 => 1,
			153 => 0,
			154 => 1,
			155 => -1,
			156 => -8,
			157 => 2,
			158 => 2,
			159 => 1,
			160 => 1,
			161 => 7,
			162 => -1,
			163 => -2,
			164 => 0,
			165 => -3,
			166 => -1,
			167 => 0,
			168 => 2,
			169 => 6,
			170 => -8,
			171 => 8,
			172 => 0,
			173 => 0,
			174 => -1,
			175 => 0,
			176 => 3,
			177 => -6,
			178 => 4,
			179 => 0,
			180 => -9,
			181 => 16,
			182 => 1,
			183 => -5,
			184 => 2,
			185 => 0,
			186 => -5,
			187 => -2,
			188 => 0,
			189 => 1,
			190 => -4,
			191 => -1,
			--Neuron 4
			192 => -2,
			193 => -6,
			194 => 15,
			195 => -1,
			196 => -14,
			197 => -5,
			198 => -8,
			199 => 8,
			200 => -6,
			201 => -2,
			202 => -4,
			203 => -3,
			204 => -2,
			205 => -2,
			206 => 0,
			207 => -12,
			208 => 17,
			209 => -2,
			210 => -2,
			211 => -4,
			212 => -7,
			213 => 4,
			214 => -6,
			215 => 4,
			216 => 0,
			217 => -2,
			218 => 0,
			219 => 5,
			220 => 10,
			221 => 4,
			222 => 3,
			223 => -1,
			224 => -1,
			225 => 10,
			226 => -3,
			227 => -4,
			228 => -1,
			229 => -5,
			230 => 4,
			231 => 3,
			232 => 0,
			233 => 9,
			234 => 9,
			235 => 3,
			236 => 4,
			237 => -2,
			238 => -1,
			239 => -1,
			240 => -4,
			241 => 4,
			242 => -1,
			243 => 2,
			244 => -1,
			245 => 6,
			246 => 0,
			247 => -5,
			248 => 1,
			249 => 0,
			250 => -6,
			251 => -1,
			252 => 0,
			253 => 0,
			254 => -1,
			255 => -1,
			--Neuron 5
			256 => 8,
			257 => 9,
			258 => 0,
			259 => -2,
			260 => -1,
			261 => -2,
			262 => -7,
			263 => 8,
			264 => 2,
			265 => -7,
			266 => 5,
			267 => 4,
			268 => -2,
			269 => 7,
			270 => 7,
			271 => 12,
			272 => -2,
			273 => 0,
			274 => -1,
			275 => -11,
			276 => -7,
			277 => -1,
			278 => 4,
			279 => 3,
			280 => -3,
			281 => -3,
			282 => 1,
			283 => 5,
			284 => -7,
			285 => 1,
			286 => 0,
			287 => 0,
			288 => 0,
			289 => 7,
			290 => 0,
			291 => 2,
			292 => -2,
			293 => -7,
			294 => -1,
			295 => 1,
			296 => 3,
			297 => 9,
			298 => -8,
			299 => 3,
			300 => -3,
			301 => -1,
			302 => 1,
			303 => 0,
			304 => 1,
			305 => -8,
			306 => 4,
			307 => 10,
			308 => 12,
			309 => -8,
			310 => 0,
			311 => 0,
			312 => 5,
			313 => 1,
			314 => -6,
			315 => 2,
			316 => 3,
			317 => 3,
			318 => 6,
			319 => 0,
			--Layer 2
			--Neuron 1
			320 => -54,
			321 => -2,
			322 => -30,
			323 => -19,
			324 => -28,
			325 => 28,
			--Neuron 2
			326 => 45,
			327 => 4,
			328 => -13,
			329 => -5,
			330 => 0,
			331 => -34,
			--Neuron 3
			332 => -20,
			333 => 16,
			334 => -43,
			335 => -23,
			336 => 31,
			337 => -23,
			--Neuron 4
			338 => -12,
			339 => 21,
			340 => 43,
			341 => -30,
			342 => -13,
			343 => -29,
			--Neuron 5
			344 => -22,
			345 => -18,
			346 => -4,
			347 => 48,
			348 => -5,
			349 => -29,
			--Neuron 6
			350 => -11,
			351 => -11,
			352 => -44,
			353 => -24,
			354 => -35,
			355 => 30);
end package NNFFPGA_Network_secondModel_statics;

-- NNFFPGA_Network_firstModel_statics.vhd
-- This is an automatically generated file containing the constants for the neural network
-- The constants are generated form a Keras Network Object via the Network-2-FPGA.py script

-- Autor: Christian Woznik
-- E-Mail: christian.woznik@posteo.de
-- This file war created on 2021-12-01
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library work;
use work.NNFPGA_pkg.all;
use work.NNFPGA_statics.all;

package NNFFPGA_Network_firstModel_statics is
	-- Layer Informations
	constant c_networkfirstModelLayerInformation : t_networkInformation(0 to 1) := (
			0 => (activationFunction => 1, inputCount => 49, neuronCount =>10),
			1 => (activationFunction => 4, inputCount => 10, neuronCount =>7));


	-- Weights Array
	constant c_networkfirstModelWeights : t_variableSizeIntegerArray(0 to 576) := (
			--Layer 1
			--Neuron 1
			0 => 6,
			1 => -1,
			2 => 1,
			3 => 10,
			4 => 5,
			5 => 0,
			6 => 6,
			7 => -2,
			8 => -18,
			9 => -5,
			10 => -2,
			11 => 4,
			12 => -8,
			13 => -1,
			14 => -4,
			15 => -14,
			16 => -18,
			17 => 6,
			18 => 5,
			19 => -17,
			20 => -2,
			21 => -16,
			22 => -35,
			23 => -31,
			24 => 2,
			25 => -2,
			26 => -31,
			27 => -7,
			28 => -9,
			29 => -22,
			30 => -19,
			31 => 6,
			32 => 4,
			33 => -24,
			34 => -5,
			35 => -5,
			36 => -13,
			37 => -16,
			38 => 1,
			39 => 2,
			40 => -10,
			41 => 2,
			42 => 1,
			43 => -5,
			44 => -1,
			45 => 3,
			46 => 7,
			47 => -3,
			48 => 1,
			49 => 65,
			--Neuron 2
			50 => -5,
			51 => -12,
			52 => 2,
			53 => 1,
			54 => 0,
			55 => -11,
			56 => -4,
			57 => -12,
			58 => -21,
			59 => 2,
			60 => -13,
			61 => 3,
			62 => -22,
			63 => -10,
			64 => -11,
			65 => -30,
			66 => 1,
			67 => -23,
			68 => -3,
			69 => -31,
			70 => -15,
			71 => 6,
			72 => -16,
			73 => 1,
			74 => -42,
			75 => -8,
			76 => -17,
			77 => 0,
			78 => -2,
			79 => -6,
			80 => 19,
			81 => 8,
			82 => 14,
			83 => -8,
			84 => -5,
			85 => -7,
			86 => -10,
			87 => 10,
			88 => 4,
			89 => 6,
			90 => -14,
			91 => -6,
			92 => 0,
			93 => -4,
			94 => 8,
			95 => 5,
			96 => 9,
			97 => -6,
			98 => -1,
			99 => 58,
			--Neuron 3
			100 => -11,
			101 => -17,
			102 => -9,
			103 => -4,
			104 => -20,
			105 => -18,
			106 => -15,
			107 => -21,
			108 => -4,
			109 => 25,
			110 => 37,
			111 => 3,
			112 => -3,
			113 => -25,
			114 => 4,
			115 => 6,
			116 => 31,
			117 => 35,
			118 => 8,
			119 => 8,
			120 => 4,
			121 => -2,
			122 => -10,
			123 => 3,
			124 => 4,
			125 => -21,
			126 => -2,
			127 => 6,
			128 => -5,
			129 => -7,
			130 => 11,
			131 => 21,
			132 => -29,
			133 => 0,
			134 => 2,
			135 => -15,
			136 => -19,
			137 => 4,
			138 => 12,
			139 => -17,
			140 => -18,
			141 => -14,
			142 => -4,
			143 => -8,
			144 => 8,
			145 => 12,
			146 => -7,
			147 => -5,
			148 => -3,
			149 => -27,
			--Neuron 4
			150 => -13,
			151 => 17,
			152 => 14,
			153 => 3,
			154 => -1,
			155 => 16,
			156 => 4,
			157 => 16,
			158 => 9,
			159 => 12,
			160 => -5,
			161 => 11,
			162 => 3,
			163 => 13,
			164 => 20,
			165 => 13,
			166 => -21,
			167 => 5,
			168 => 3,
			169 => 4,
			170 => 2,
			171 => -5,
			172 => 4,
			173 => -3,
			174 => -14,
			175 => -2,
			176 => -5,
			177 => -3,
			178 => 0,
			179 => -1,
			180 => -1,
			181 => 2,
			182 => -21,
			183 => 16,
			184 => 9,
			185 => 12,
			186 => 1,
			187 => 5,
			188 => 7,
			189 => 11,
			190 => 10,
			191 => 13,
			192 => 19,
			193 => 17,
			194 => 0,
			195 => 2,
			196 => 26,
			197 => 17,
			198 => -14,
			199 => -60,
			--Neuron 5
			200 => 16,
			201 => 10,
			202 => 23,
			203 => 4,
			204 => 20,
			205 => 1,
			206 => 14,
			207 => 16,
			208 => 13,
			209 => 3,
			210 => 1,
			211 => -24,
			212 => 13,
			213 => 14,
			214 => -11,
			215 => 6,
			216 => 16,
			217 => 4,
			218 => -12,
			219 => 0,
			220 => -12,
			221 => -25,
			222 => -24,
			223 => -12,
			224 => 9,
			225 => -41,
			226 => -27,
			227 => -32,
			228 => -15,
			229 => -2,
			230 => 12,
			231 => 27,
			232 => -9,
			233 => -17,
			234 => -17,
			235 => -6,
			236 => 10,
			237 => 14,
			238 => 6,
			239 => 2,
			240 => -2,
			241 => -3,
			242 => 5,
			243 => 13,
			244 => 24,
			245 => 9,
			246 => 8,
			247 => 5,
			248 => 17,
			249 => 12,
			--Neuron 6
			250 => -13,
			251 => -19,
			252 => -8,
			253 => -7,
			254 => -12,
			255 => -19,
			256 => -13,
			257 => 1,
			258 => 5,
			259 => -8,
			260 => -10,
			261 => -9,
			262 => 6,
			263 => 1,
			264 => 14,
			265 => 16,
			266 => 2,
			267 => -8,
			268 => 3,
			269 => 18,
			270 => 16,
			271 => 10,
			272 => 15,
			273 => 14,
			274 => 12,
			275 => 14,
			276 => 13,
			277 => 12,
			278 => 1,
			279 => 4,
			280 => -2,
			281 => 11,
			282 => 1,
			283 => 6,
			284 => -3,
			285 => -3,
			286 => -17,
			287 => -23,
			288 => -25,
			289 => -26,
			290 => -15,
			291 => -6,
			292 => -11,
			293 => -18,
			294 => -10,
			295 => -5,
			296 => -12,
			297 => -18,
			298 => -15,
			299 => 2,
			--Neuron 7
			300 => 11,
			301 => -15,
			302 => -5,
			303 => -9,
			304 => -3,
			305 => -14,
			306 => 10,
			307 => -15,
			308 => 20,
			309 => 18,
			310 => 27,
			311 => 18,
			312 => 23,
			313 => -12,
			314 => 1,
			315 => 7,
			316 => -6,
			317 => -22,
			318 => -6,
			319 => 9,
			320 => 2,
			321 => 5,
			322 => 8,
			323 => -10,
			324 => 23,
			325 => -6,
			326 => 14,
			327 => 4,
			328 => 9,
			329 => -5,
			330 => 9,
			331 => -25,
			332 => 9,
			333 => -5,
			334 => 17,
			335 => -6,
			336 => 25,
			337 => -8,
			338 => 2,
			339 => -14,
			340 => 21,
			341 => -4,
			342 => 4,
			343 => -18,
			344 => 0,
			345 => -4,
			346 => -2,
			347 => -13,
			348 => 12,
			349 => -47,
			--Neuron 8
			350 => 7,
			351 => 0,
			352 => 3,
			353 => 7,
			354 => 5,
			355 => -3,
			356 => 9,
			357 => 4,
			358 => 7,
			359 => -2,
			360 => 4,
			361 => -4,
			362 => 5,
			363 => 5,
			364 => 11,
			365 => 12,
			366 => -11,
			367 => -4,
			368 => -15,
			369 => 12,
			370 => 6,
			371 => 8,
			372 => 3,
			373 => -23,
			374 => -61,
			375 => -31,
			376 => 2,
			377 => 3,
			378 => 3,
			379 => -3,
			380 => -30,
			381 => -32,
			382 => -31,
			383 => -3,
			384 => 1,
			385 => -3,
			386 => -3,
			387 => -17,
			388 => -13,
			389 => -17,
			390 => -2,
			391 => -4,
			392 => 5,
			393 => -1,
			394 => 6,
			395 => 18,
			396 => 12,
			397 => -1,
			398 => 0,
			399 => 58,
			--Neuron 9
			400 => 0,
			401 => -4,
			402 => 6,
			403 => -8,
			404 => 7,
			405 => 0,
			406 => 0,
			407 => -6,
			408 => -18,
			409 => 1,
			410 => -13,
			411 => 13,
			412 => -15,
			413 => -14,
			414 => -24,
			415 => -12,
			416 => 27,
			417 => 12,
			418 => 21,
			419 => -12,
			420 => -6,
			421 => -5,
			422 => -2,
			423 => 23,
			424 => -14,
			425 => 18,
			426 => -21,
			427 => -12,
			428 => 12,
			429 => 8,
			430 => 7,
			431 => -29,
			432 => 22,
			433 => 1,
			434 => -10,
			435 => 16,
			436 => -15,
			437 => 5,
			438 => -26,
			439 => 5,
			440 => 3,
			441 => 5,
			442 => -8,
			443 => -5,
			444 => 1,
			445 => -13,
			446 => 4,
			447 => -8,
			448 => -15,
			449 => 1,
			--Neuron 10
			450 => 3,
			451 => 4,
			452 => 12,
			453 => 12,
			454 => 12,
			455 => 3,
			456 => 0,
			457 => -3,
			458 => -9,
			459 => -4,
			460 => -3,
			461 => 10,
			462 => 8,
			463 => 2,
			464 => -6,
			465 => 4,
			466 => -12,
			467 => -21,
			468 => -26,
			469 => 6,
			470 => 8,
			471 => 6,
			472 => 19,
			473 => -24,
			474 => -29,
			475 => -22,
			476 => 2,
			477 => 8,
			478 => 17,
			479 => 18,
			480 => 2,
			481 => -12,
			482 => 2,
			483 => 4,
			484 => 17,
			485 => 6,
			486 => 20,
			487 => 21,
			488 => 26,
			489 => 23,
			490 => 4,
			491 => 11,
			492 => -11,
			493 => 3,
			494 => 9,
			495 => 6,
			496 => -9,
			497 => 2,
			498 => 10,
			499 => -45,
			--Layer 2
			--Neuron 1
			500 => -61,
			501 => -62,
			502 => -47,
			503 => -43,
			504 => -52,
			505 => -57,
			506 => -57,
			507 => -34,
			508 => -72,
			509 => -60,
			510 => -113,
			--Neuron 2
			511 => -114,
			512 => -93,
			513 => -9,
			514 => 38,
			515 => -2,
			516 => -113,
			517 => 20,
			518 => 33,
			519 => -71,
			520 => 61,
			521 => -63,
			--Neuron 3
			522 => -53,
			523 => -117,
			524 => -85,
			525 => 43,
			526 => 21,
			527 => -120,
			528 => 29,
			529 => -88,
			530 => 6,
			531 => -108,
			532 => 17,
			--Neuron 4
			533 => -68,
			534 => -92,
			535 => 40,
			536 => -111,
			537 => -116,
			538 => -20,
			539 => 20,
			540 => 15,
			541 => 29,
			542 => -77,
			543 => 37,
			--Neuron 5
			544 => -81,
			545 => 15,
			546 => -77,
			547 => -68,
			548 => -38,
			549 => 35,
			550 => -51,
			551 => -51,
			552 => -81,
			553 => 26,
			554 => 48,
			--Neuron 6
			555 => 32,
			556 => 21,
			557 => 48,
			558 => -71,
			559 => 13,
			560 => -77,
			561 => -74,
			562 => -83,
			563 => 29,
			564 => -87,
			565 => -34,
			--Neuron 7
			566 => 38,
			567 => 3,
			568 => -79,
			569 => -62,
			570 => 1,
			571 => -36,
			572 => -55,
			573 => 27,
			574 => -24,
			575 => -46,
			576 => 58);
end package NNFFPGA_Network_firstModel_statics;
